magic
tech sky130A
magscale 1 2
timestamp 1747152884
<< error_p >>
rect -29 -211 29 -205
rect -29 -245 -17 -211
rect -29 -251 29 -245
<< nwell >>
rect -211 -384 211 384
<< pmoshvt >>
rect -15 -164 15 236
<< pdiff >>
rect -73 224 -15 236
rect -73 -152 -61 224
rect -27 -152 -15 224
rect -73 -164 -15 -152
rect 15 224 73 236
rect 15 -152 27 224
rect 61 -152 73 224
rect 15 -164 73 -152
<< pdiffc >>
rect -61 -152 -27 224
rect 27 -152 61 224
<< nsubdiff >>
rect -175 314 -79 348
rect 79 314 175 348
rect -175 251 -141 314
rect 141 251 175 314
rect -175 -314 -141 -251
rect 141 -314 175 -251
rect -175 -348 -79 -314
rect 79 -348 175 -314
<< nsubdiffcont >>
rect -79 314 79 348
rect -175 -251 -141 251
rect 141 -251 175 251
rect -79 -348 79 -314
<< poly >>
rect -15 236 15 262
rect -15 -195 15 -164
rect -33 -211 33 -195
rect -33 -245 -17 -211
rect 17 -245 33 -211
rect -33 -261 33 -245
<< polycont >>
rect -17 -245 17 -211
<< locali >>
rect -175 314 -79 348
rect 79 314 175 348
rect -175 251 -141 314
rect 141 251 175 314
rect -61 224 -27 240
rect -61 -168 -27 -152
rect 27 224 61 240
rect 27 -168 61 -152
rect -33 -245 -17 -211
rect 17 -245 33 -211
rect -175 -314 -141 -251
rect 141 -314 175 -251
rect -175 -348 -79 -314
rect 79 -348 175 -314
<< viali >>
rect -61 -152 -27 224
rect 27 -152 61 224
rect -17 -245 17 -211
<< metal1 >>
rect -67 224 -21 236
rect -67 -152 -61 224
rect -27 -152 -21 224
rect -67 -164 -21 -152
rect 21 224 67 236
rect 21 -152 27 224
rect 61 -152 67 224
rect 21 -164 67 -152
rect -29 -211 29 -205
rect -29 -245 -17 -211
rect 17 -245 29 -211
rect -29 -251 29 -245
<< properties >>
string FIXED_BBOX -158 -331 158 331
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 2.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
